module COMPARE (lt, gt, eq, data1, data2);
  
